module LEG(
	input i_clk
);
endmodule
